magic
tech scmos
timestamp 1571845397
<< nwell >>
rect -4 34 38 68
<< pwell >>
rect -4 68 38 132
rect -4 0 38 34
<< ntransistor >>
rect 16 105 18 109
rect 24 105 26 109
rect 16 77 18 81
rect 24 77 26 81
rect 16 24 18 28
<< ptransistor >>
rect 8 56 10 60
rect 16 56 18 60
rect 24 56 26 60
rect 16 40 18 44
<< ndiffusion >>
rect 15 105 16 109
rect 18 105 19 109
rect 23 105 24 109
rect 26 105 27 109
rect 15 77 16 81
rect 18 77 19 81
rect 23 77 24 81
rect 26 80 31 81
rect 26 77 27 80
rect 15 24 16 28
rect 18 24 19 28
<< pdiffusion >>
rect 7 56 8 60
rect 10 56 11 60
rect 15 56 16 60
rect 18 56 19 60
rect 23 56 24 60
rect 26 56 27 60
rect 15 40 16 44
rect 18 40 19 44
<< ndcontact >>
rect 11 105 15 109
rect 19 105 23 109
rect 27 105 31 109
rect 11 77 15 81
rect 19 77 23 81
rect 27 76 31 80
rect 11 24 15 28
rect 19 24 23 28
<< pdcontact >>
rect 3 56 7 60
rect 11 56 15 60
rect 19 56 23 60
rect 27 56 31 60
rect 11 40 15 44
rect 19 40 23 44
<< psubstratepcontact >>
rect 8 120 12 124
rect 3 18 7 22
<< nsubstratencontact >>
rect 27 48 31 52
<< polysilicon >>
rect 16 109 18 111
rect 24 109 26 112
rect 16 102 18 105
rect 24 103 26 105
rect 16 81 18 84
rect 24 81 26 83
rect 8 60 10 62
rect 16 60 18 77
rect 24 70 26 77
rect 24 66 25 70
rect 24 60 26 66
rect 8 36 10 56
rect 16 54 18 56
rect 24 54 26 56
rect 16 44 18 46
rect 16 28 18 40
rect 16 14 18 24
<< polycontact >>
rect 23 112 27 116
rect 15 98 19 102
rect 15 84 19 88
rect 25 66 29 70
rect 8 32 12 36
rect 15 10 19 14
<< metal1 >>
rect 0 121 4 124
rect 12 121 34 124
rect 12 120 14 121
rect 11 109 14 120
rect 0 95 34 98
rect 0 88 34 90
rect 0 87 15 88
rect 19 87 34 88
rect 0 67 25 70
rect 29 67 34 70
rect 3 52 6 56
rect 27 52 31 56
rect 0 48 27 52
rect 31 48 34 52
rect 19 44 23 48
rect 11 36 14 40
rect 12 32 14 36
rect 11 28 14 32
rect 19 21 22 24
rect 7 18 22 21
rect 0 11 15 14
rect 19 11 34 14
<< m2contact >>
rect 4 120 8 124
rect 19 112 23 116
rect 27 101 31 105
rect 27 80 31 84
rect 11 73 15 77
rect 11 60 15 64
rect 3 22 7 26
<< metal2 >>
rect 27 127 31 132
rect 4 26 7 120
rect 27 116 31 123
rect 23 112 31 116
rect 28 84 31 101
rect 11 64 14 73
rect 11 51 14 60
rect 11 48 29 51
rect 26 0 29 48
<< m3contact >>
rect 27 123 31 127
<< metal3 >>
rect 26 127 32 132
rect 26 123 27 127
rect 31 123 32 127
rect 26 122 32 123
<< m3p >>
rect 0 0 34 132
<< labels >>
rlabel metal1 34 11 34 11 8 reset
rlabel metal2 29 0 29 0 1 Q
rlabel metal1 34 67 34 67 7 en2_M
rlabel metal1 34 95 34 95 7 M
rlabel metal1 34 121 34 121 5 gnd
rlabel metal1 34 48 34 48 5 vdd
rlabel metal1 34 87 34 87 7 en1_M
rlabel metal2 31 132 31 132 5 D
<< end >>
