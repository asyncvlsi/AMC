magic
tech scmos
timestamp 1561575115
<< nwell >>
rect 0 116 66 160
rect 0 24 66 68
<< pwell >>
rect 0 160 66 186
rect 0 68 66 116
rect 0 -2 66 24
<< ntransistor >>
rect 15 171 17 179
rect 23 171 25 179
rect 39 175 41 179
rect 47 175 49 179
rect 15 97 17 105
rect 23 97 25 105
rect 39 97 41 101
rect 47 97 49 101
rect 15 79 17 87
rect 23 79 25 87
rect 39 83 41 87
rect 47 83 49 87
rect 15 5 17 13
rect 23 5 25 13
rect 39 5 41 9
rect 47 5 49 9
<< ptransistor >>
rect 15 143 17 151
rect 23 143 25 151
rect 39 143 41 151
rect 47 143 49 151
rect 15 125 17 133
rect 23 125 25 133
rect 39 125 41 133
rect 47 125 49 133
rect 15 51 17 59
rect 23 51 25 59
rect 39 51 41 59
rect 47 51 49 59
rect 15 33 17 41
rect 23 33 25 41
rect 39 33 41 41
rect 47 33 49 41
<< ndiffusion >>
rect 10 177 15 179
rect 14 173 15 177
rect 10 171 15 173
rect 17 177 23 179
rect 17 173 18 177
rect 22 173 23 177
rect 17 171 23 173
rect 25 177 30 179
rect 25 173 26 177
rect 38 175 39 179
rect 41 175 42 179
rect 46 175 47 179
rect 49 175 50 179
rect 25 171 30 173
rect 10 103 15 105
rect 14 99 15 103
rect 10 97 15 99
rect 17 103 23 105
rect 17 99 18 103
rect 22 99 23 103
rect 17 97 23 99
rect 25 103 30 105
rect 25 99 26 103
rect 25 97 30 99
rect 38 97 39 101
rect 41 97 42 101
rect 46 97 47 101
rect 49 97 50 101
rect 14 79 15 87
rect 17 85 23 87
rect 17 81 18 85
rect 22 81 23 85
rect 17 79 23 81
rect 25 85 30 87
rect 25 81 26 85
rect 38 83 39 87
rect 41 83 42 87
rect 46 83 47 87
rect 49 83 50 87
rect 25 79 30 81
rect 10 11 15 13
rect 14 7 15 11
rect 10 5 15 7
rect 17 11 23 13
rect 17 7 18 11
rect 22 7 23 11
rect 17 5 23 7
rect 25 11 30 13
rect 25 7 26 11
rect 25 5 30 7
rect 38 5 39 9
rect 41 5 42 9
rect 46 5 47 9
rect 49 5 50 9
<< pdiffusion >>
rect 10 149 15 151
rect 14 145 15 149
rect 10 143 15 145
rect 17 149 23 151
rect 17 145 18 149
rect 22 145 23 149
rect 17 143 23 145
rect 25 149 30 151
rect 25 145 26 149
rect 25 143 30 145
rect 34 149 39 151
rect 38 145 39 149
rect 34 143 39 145
rect 41 149 47 151
rect 41 145 42 149
rect 46 145 47 149
rect 41 143 47 145
rect 49 149 54 151
rect 49 145 50 149
rect 49 143 54 145
rect 10 131 15 133
rect 14 127 15 131
rect 10 125 15 127
rect 17 131 23 133
rect 17 127 18 131
rect 22 127 23 131
rect 17 125 23 127
rect 25 131 30 133
rect 25 127 26 131
rect 25 125 30 127
rect 34 131 39 133
rect 38 127 39 131
rect 34 125 39 127
rect 41 131 47 133
rect 41 127 42 131
rect 46 127 47 131
rect 41 125 47 127
rect 49 131 54 133
rect 49 127 50 131
rect 49 125 54 127
rect 10 55 15 59
rect 14 51 15 55
rect 17 57 23 59
rect 17 53 18 57
rect 22 53 23 57
rect 17 51 23 53
rect 25 57 30 59
rect 25 53 26 57
rect 25 51 30 53
rect 34 57 39 59
rect 38 53 39 57
rect 34 51 39 53
rect 41 57 47 59
rect 41 53 42 57
rect 46 53 47 57
rect 41 51 47 53
rect 49 57 54 59
rect 49 53 50 57
rect 49 51 54 53
rect 10 39 15 41
rect 14 35 15 39
rect 10 33 15 35
rect 17 39 23 41
rect 17 35 18 39
rect 22 35 23 39
rect 17 33 23 35
rect 25 39 30 41
rect 25 35 26 39
rect 25 33 30 35
rect 34 39 39 41
rect 38 35 39 39
rect 34 33 39 35
rect 41 39 47 41
rect 41 35 42 39
rect 46 35 47 39
rect 41 33 47 35
rect 49 39 54 41
rect 49 35 50 39
rect 49 33 54 35
<< ndcontact >>
rect 10 173 14 177
rect 18 173 22 177
rect 26 173 30 177
rect 34 175 38 179
rect 42 175 46 179
rect 50 175 54 179
rect 10 99 14 103
rect 18 99 22 103
rect 26 99 30 103
rect 34 97 38 101
rect 42 97 46 101
rect 50 97 54 101
rect 10 79 14 87
rect 18 81 22 85
rect 26 81 30 85
rect 34 83 38 87
rect 42 83 46 87
rect 50 83 54 87
rect 10 7 14 11
rect 18 7 22 11
rect 26 7 30 11
rect 34 5 38 9
rect 42 5 46 9
rect 50 5 54 9
<< pdcontact >>
rect 10 145 14 149
rect 18 145 22 149
rect 26 145 30 149
rect 34 145 38 149
rect 42 145 46 149
rect 50 145 54 149
rect 10 127 14 131
rect 18 127 22 131
rect 26 127 30 131
rect 34 127 38 131
rect 42 127 46 131
rect 50 127 54 131
rect 10 51 14 55
rect 18 53 22 57
rect 26 53 30 57
rect 34 53 38 57
rect 42 53 46 57
rect 50 53 54 57
rect 10 35 14 39
rect 18 35 22 39
rect 26 35 30 39
rect 34 35 38 39
rect 42 35 46 39
rect 50 35 54 39
<< psubstratepcontact >>
rect 34 167 38 171
rect 34 105 38 109
rect 34 75 38 79
rect 34 13 38 17
<< nsubstratencontact >>
rect 58 145 62 149
rect 58 127 62 131
rect 58 53 62 57
rect 58 35 62 39
<< polysilicon >>
rect 15 179 17 181
rect 23 179 25 181
rect 39 179 41 181
rect 47 179 49 181
rect 15 151 17 171
rect 23 166 25 171
rect 24 162 25 166
rect 23 151 25 162
rect 39 162 41 175
rect 47 162 49 175
rect 39 160 49 162
rect 39 151 41 160
rect 47 151 49 160
rect 15 141 17 143
rect 23 141 25 143
rect 39 141 41 143
rect 47 141 49 143
rect 15 133 17 135
rect 23 133 25 135
rect 39 133 41 135
rect 47 133 49 135
rect 15 105 17 125
rect 23 114 25 125
rect 24 110 25 114
rect 39 116 41 125
rect 47 116 49 125
rect 39 114 49 116
rect 23 105 25 110
rect 39 101 41 114
rect 47 101 49 114
rect 15 95 17 97
rect 23 95 25 97
rect 39 95 41 97
rect 47 95 49 97
rect 15 87 17 89
rect 23 87 25 89
rect 39 87 41 89
rect 47 87 49 89
rect 15 59 17 79
rect 23 76 25 79
rect 24 72 25 76
rect 23 59 25 72
rect 39 70 41 83
rect 47 70 49 83
rect 39 68 49 70
rect 39 59 41 68
rect 47 59 49 68
rect 15 49 17 51
rect 23 49 25 51
rect 39 49 41 51
rect 47 49 49 51
rect 15 41 17 43
rect 23 41 25 43
rect 39 41 41 43
rect 47 41 49 43
rect 15 13 17 33
rect 23 22 25 33
rect 24 18 25 22
rect 39 24 41 33
rect 47 24 49 33
rect 39 22 49 24
rect 23 13 25 18
rect 39 9 41 22
rect 47 9 49 22
rect 15 3 17 5
rect 23 3 25 5
rect 39 3 41 5
rect 47 3 49 5
<< polycontact >>
rect 11 154 15 158
rect 20 162 24 166
rect 35 159 39 163
rect 11 118 15 122
rect 20 110 24 114
rect 35 113 39 117
rect 11 62 15 66
rect 20 72 24 76
rect 35 67 39 71
rect 11 26 15 30
rect 20 18 24 22
rect 35 21 39 25
<< metal1 >>
rect 0 182 66 186
rect 10 177 14 182
rect 34 179 38 182
rect 50 179 54 182
rect 4 162 20 165
rect 27 162 30 173
rect 34 171 38 175
rect 57 175 66 179
rect 42 170 46 175
rect 57 170 61 175
rect 42 167 61 170
rect 27 159 35 162
rect 27 157 30 159
rect 18 154 30 157
rect 18 149 22 154
rect 34 149 38 151
rect 10 140 14 145
rect 26 140 30 145
rect 34 140 38 145
rect 42 149 46 167
rect 42 143 46 145
rect 50 140 54 145
rect 58 140 62 145
rect 0 136 66 140
rect 10 131 14 136
rect 26 131 30 136
rect 34 131 38 136
rect 18 122 22 127
rect 34 125 38 127
rect 42 131 46 133
rect 50 131 54 136
rect 58 131 62 136
rect 18 119 30 122
rect 27 117 30 119
rect 27 114 35 117
rect 4 110 20 113
rect 27 103 30 114
rect 42 109 46 127
rect 34 101 38 105
rect 10 94 14 99
rect 42 106 61 109
rect 42 101 46 106
rect 57 101 61 106
rect 57 97 66 101
rect 34 94 38 97
rect 50 94 54 97
rect 0 90 66 94
rect 10 87 14 90
rect 34 87 38 90
rect 50 87 54 90
rect 4 73 20 76
rect 27 70 30 81
rect 34 79 38 83
rect 57 83 66 87
rect 42 78 46 83
rect 57 78 61 83
rect 42 75 61 78
rect 0 65 11 68
rect 27 67 35 70
rect 27 65 30 67
rect 18 62 30 65
rect 18 57 22 62
rect 34 57 38 59
rect 10 48 14 51
rect 26 48 30 53
rect 34 48 38 53
rect 42 57 46 75
rect 42 51 46 53
rect 50 48 54 53
rect 58 48 62 53
rect 0 44 66 48
rect 10 39 14 44
rect 26 39 30 44
rect 34 39 38 44
rect 18 30 22 35
rect 34 33 38 35
rect 42 39 46 41
rect 50 39 54 44
rect 58 39 62 44
rect 18 27 30 30
rect 27 25 30 27
rect 27 22 35 25
rect 4 19 20 22
rect 27 11 30 22
rect 42 17 46 35
rect 34 9 38 13
rect 10 2 14 7
rect 42 14 60 17
rect 42 9 46 14
rect 57 9 60 14
rect 57 5 66 9
rect 34 2 38 5
rect 50 2 54 5
rect 0 -2 66 2
<< m2contact >>
rect 0 162 4 166
rect 7 154 11 158
rect 7 118 11 122
rect 0 110 4 114
rect 0 73 4 77
rect 11 66 15 70
rect 7 26 11 30
rect 0 19 4 23
<< metal2 >>
rect 11 70 15 158
rect 11 26 15 66
<< m3contact >>
rect 4 162 8 166
rect 4 110 8 114
rect 4 73 8 77
rect 4 19 8 23
<< metal3 >>
rect 0 166 9 167
rect 0 162 4 166
rect 8 162 9 166
rect 0 161 9 162
rect 0 114 9 115
rect 0 110 4 114
rect 8 110 9 114
rect 0 109 9 110
rect 0 77 9 78
rect 0 73 4 77
rect 8 73 9 77
rect 0 72 9 73
rect 0 23 9 24
rect 0 19 4 23
rect 8 19 9 23
rect 0 18 9 19
<< m3p >>
rect 0 0 66 184
<< labels >>
rlabel m2contact 0 162 0 162 3 in3
rlabel metal1 0 184 0 184 2 gnd
rlabel metal1 0 138 0 138 2 vdd
rlabel m2contact 0 110 0 110 3 in2
rlabel metal1 0 46 0 46 2 vdd
rlabel m2contact 0 19 0 19 3 in0
rlabel metal1 0 0 0 0 6 gnd
rlabel metal1 0 92 0 92 4 gnd
rlabel m2contact 0 73 0 73 3 in1
rlabel metal1 0 65 0 65 3 en
rlabel metal1 66 175 66 175 7 out3
rlabel metal1 66 84 66 84 1 out1
rlabel metal1 66 97 66 97 7 out2
rlabel metal1 66 5 66 5 7 out0
<< end >>
