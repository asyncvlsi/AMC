magic
tech scmos
timestamp 1564444365
<< nwell >>
rect -6 107 34 252
rect -6 30 34 62
<< pwell >>
rect -6 252 34 309
rect -6 62 34 107
rect -6 0 34 30
<< ntransistor >>
rect 12 280 14 298
rect 12 258 14 267
rect 20 258 22 267
rect 9 97 11 101
rect 17 97 19 101
rect 13 16 15 24
rect 21 16 23 24
<< ptransistor >>
rect 12 228 14 246
rect 20 228 22 246
rect 10 178 12 202
rect 21 147 23 171
rect 9 113 11 121
rect 17 113 19 121
rect 13 36 15 44
rect 21 36 23 44
<< ndiffusion >>
rect 11 280 12 298
rect 14 280 15 298
rect 11 258 12 267
rect 14 258 15 267
rect 19 258 20 267
rect 22 258 23 267
rect 8 97 9 101
rect 11 97 12 101
rect 16 97 17 101
rect 19 97 20 101
rect 12 16 13 24
rect 15 16 16 24
rect 20 16 21 24
rect 23 16 24 24
<< pdiffusion >>
rect 7 244 12 246
rect 11 230 12 244
rect 7 228 12 230
rect 14 244 20 246
rect 14 230 15 244
rect 19 230 20 244
rect 14 228 20 230
rect 22 244 27 246
rect 22 230 23 244
rect 22 228 27 230
rect 9 178 10 202
rect 12 178 13 202
rect 20 147 21 171
rect 23 147 24 171
rect 8 113 9 121
rect 11 113 12 121
rect 16 113 17 121
rect 19 113 20 121
rect 8 42 13 44
rect 12 38 13 42
rect 8 36 13 38
rect 15 42 21 44
rect 15 38 16 42
rect 20 38 21 42
rect 15 36 21 38
rect 23 42 28 44
rect 23 38 24 42
rect 23 36 28 38
<< ndcontact >>
rect 7 280 11 298
rect 15 280 19 298
rect 7 258 11 267
rect 15 258 19 267
rect 23 258 27 267
rect 4 97 8 101
rect 12 97 16 101
rect 20 97 24 101
rect 8 16 12 24
rect 16 16 20 24
rect 24 16 28 24
<< pdcontact >>
rect 7 230 11 244
rect 15 230 19 244
rect 23 230 27 244
rect 5 178 9 202
rect 13 178 17 202
rect 16 147 20 171
rect 24 147 28 171
rect 4 113 8 121
rect 12 113 16 121
rect 20 113 24 121
rect 8 38 12 42
rect 16 38 20 42
rect 24 38 28 42
<< psubstratepcontact >>
rect -2 297 2 301
rect 16 83 20 87
rect -2 16 2 20
<< nsubstratencontact >>
rect 12 212 16 216
rect 12 135 16 139
rect 27 48 31 52
<< polysilicon >>
rect 12 298 14 300
rect 12 279 14 280
rect 12 277 31 279
rect 3 272 22 274
rect 3 255 5 272
rect 12 267 14 269
rect 20 267 22 272
rect 3 251 4 255
rect 3 209 5 251
rect 12 246 14 258
rect 20 246 22 258
rect 12 223 14 228
rect 20 226 22 228
rect 12 221 22 223
rect 23 205 25 219
rect 10 202 12 204
rect 10 146 12 178
rect 29 174 31 277
rect 21 172 31 174
rect 21 171 23 172
rect 21 146 23 147
rect 10 144 27 146
rect 5 128 7 139
rect 25 132 27 144
rect 5 126 31 128
rect 9 121 11 123
rect 17 121 19 123
rect 9 101 11 113
rect 17 110 19 113
rect 18 106 19 110
rect 17 101 19 106
rect 4 79 6 90
rect 4 64 6 75
rect 9 71 11 97
rect 17 95 19 97
rect 4 62 15 64
rect 29 62 31 126
rect 13 44 15 58
rect 21 58 27 60
rect 21 44 23 58
rect 13 34 15 36
rect 6 28 15 30
rect 13 24 15 28
rect 21 24 23 36
rect 13 14 15 16
rect 21 9 23 16
rect 7 7 23 9
<< polycontact >>
rect 4 251 8 255
rect 22 219 26 223
rect 3 205 7 209
rect 21 201 25 205
rect 3 139 7 143
rect 21 132 25 136
rect 14 106 18 110
rect 2 90 6 94
rect 2 75 6 79
rect 9 67 13 71
rect 11 58 15 62
rect 27 58 31 62
rect 2 28 6 32
rect 3 7 7 11
<< metal1 >>
rect 2 301 34 305
rect 7 298 11 301
rect 15 267 18 280
rect 7 255 11 258
rect 8 251 11 255
rect 7 244 11 251
rect 7 228 11 230
rect 15 244 19 246
rect 23 244 27 258
rect 15 225 18 230
rect 13 222 18 225
rect 23 223 27 230
rect 13 216 16 222
rect 26 219 27 223
rect 0 212 12 216
rect 16 212 27 216
rect 31 212 34 216
rect 3 202 7 205
rect 3 178 5 202
rect 3 143 6 178
rect 25 171 28 204
rect 12 139 27 143
rect 12 121 16 135
rect 21 121 24 132
rect 4 110 8 113
rect 4 106 14 110
rect 4 101 8 106
rect 21 101 24 113
rect 4 94 8 97
rect 6 90 8 94
rect 12 87 16 97
rect 2 83 16 87
rect -2 67 9 70
rect 13 67 34 70
rect 2 32 5 67
rect 25 44 27 48
rect 25 42 28 44
rect 9 24 12 38
rect 16 24 20 38
rect 25 24 27 27
rect 12 16 13 24
rect 9 15 13 16
rect 10 11 13 15
rect 10 7 27 11
<< m2contact >>
rect -2 301 2 305
rect 27 212 31 216
rect 13 202 17 206
rect 17 171 21 175
rect 27 139 31 143
rect -2 83 2 87
rect 27 44 31 48
rect 27 24 31 28
rect -2 20 2 24
rect 27 7 31 11
rect 3 3 7 7
<< metal2 >>
rect -2 305 2 309
rect -2 87 2 301
rect -2 24 2 83
rect -2 16 2 20
rect 10 206 14 309
rect 10 202 13 206
rect -2 12 -1 16
rect 3 0 7 3
rect 10 0 14 202
rect 20 175 24 309
rect 21 171 24 175
rect 20 0 24 171
rect 27 216 31 309
rect 27 143 31 212
rect 27 48 31 139
rect 27 5 31 7
<< m3contact >>
rect -1 12 3 16
rect 27 28 31 32
rect 27 1 31 5
<< metal3 >>
rect 26 32 32 33
rect 26 28 27 32
rect 31 28 32 32
rect 26 17 32 28
rect -2 16 32 17
rect -2 12 -1 16
rect 3 12 32 16
rect -2 11 32 12
rect 26 5 32 6
rect 26 1 27 5
rect 31 1 32 5
rect 26 0 32 1
<< m3p >>
rect 0 0 34 309
<< labels >>
flabel metal1 34 212 34 212 6 FreeSans 26 180 0 0 vdd
flabel metal1 34 301 34 301 6 FreeSans 26 180 0 0 gnd
flabel metal1 34 67 34 67 6 FreeSans 26 180 0 0 en
rlabel metal3 31 0 31 0 8 dout
rlabel metal2 24 0 24 0 1 bl
rlabel metal2 7 0 7 0 1 dout_bar
rlabel metal2 13 0 13 0 1 br
<< properties >>
string path 270.000 468.000 270.000 486.000 288.000 486.000 288.000 468.000 270.000 468.000 
<< end >>
