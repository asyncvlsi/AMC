magic
tech scmos
timestamp 1551900896
<< nwell >>
rect 0 116 64 160
rect 0 24 64 68
<< pwell >>
rect 0 160 64 186
rect 0 68 64 116
rect 0 -4 64 24
<< ntransistor >>
rect 21 171 23 179
rect 29 171 31 179
rect 45 175 47 179
rect 21 97 23 105
rect 29 97 31 105
rect 45 97 47 101
rect 12 83 14 87
rect 21 79 23 87
rect 29 79 31 87
rect 45 83 47 87
rect 21 5 23 13
rect 29 5 31 13
rect 45 5 47 9
<< ptransistor >>
rect 21 143 23 151
rect 29 143 31 151
rect 45 143 47 151
rect 21 125 23 133
rect 29 125 31 133
rect 45 125 47 133
rect 12 51 14 59
rect 21 51 23 59
rect 29 51 31 59
rect 45 51 47 59
rect 21 33 23 41
rect 29 33 31 41
rect 45 33 47 41
<< ndiffusion >>
rect 16 177 21 179
rect 20 173 21 177
rect 16 171 21 173
rect 23 177 29 179
rect 23 173 24 177
rect 28 173 29 177
rect 23 171 29 173
rect 31 177 36 179
rect 31 173 32 177
rect 44 175 45 179
rect 47 175 48 179
rect 31 171 36 173
rect 16 103 21 105
rect 20 99 21 103
rect 16 97 21 99
rect 23 103 29 105
rect 23 99 24 103
rect 28 99 29 103
rect 23 97 29 99
rect 31 103 36 105
rect 31 99 32 103
rect 31 97 36 99
rect 44 97 45 101
rect 47 97 48 101
rect 11 83 12 87
rect 14 83 16 87
rect 20 79 21 87
rect 23 85 29 87
rect 23 81 24 85
rect 28 81 29 85
rect 23 79 29 81
rect 31 85 36 87
rect 31 81 32 85
rect 44 83 45 87
rect 47 83 48 87
rect 31 79 36 81
rect 16 11 21 13
rect 20 7 21 11
rect 16 5 21 7
rect 23 11 29 13
rect 23 7 24 11
rect 28 7 29 11
rect 23 5 29 7
rect 31 11 36 13
rect 31 7 32 11
rect 31 5 36 7
rect 44 5 45 9
rect 47 5 48 9
<< pdiffusion >>
rect 16 149 21 151
rect 20 145 21 149
rect 16 143 21 145
rect 23 149 29 151
rect 23 145 24 149
rect 28 145 29 149
rect 23 143 29 145
rect 31 149 36 151
rect 31 145 32 149
rect 31 143 36 145
rect 40 149 45 151
rect 44 145 45 149
rect 40 143 45 145
rect 47 149 52 151
rect 47 145 48 149
rect 47 143 52 145
rect 16 131 21 133
rect 20 127 21 131
rect 16 125 21 127
rect 23 131 29 133
rect 23 127 24 131
rect 28 127 29 131
rect 23 125 29 127
rect 31 131 36 133
rect 31 127 32 131
rect 31 125 36 127
rect 40 131 45 133
rect 44 127 45 131
rect 40 125 45 127
rect 47 131 52 133
rect 47 127 48 131
rect 47 125 52 127
rect 7 55 12 59
rect 11 51 12 55
rect 14 55 21 59
rect 14 51 16 55
rect 20 51 21 55
rect 23 57 29 59
rect 23 53 24 57
rect 28 53 29 57
rect 23 51 29 53
rect 31 57 36 59
rect 31 53 32 57
rect 31 51 36 53
rect 40 57 45 59
rect 44 53 45 57
rect 40 51 45 53
rect 47 57 52 59
rect 47 53 48 57
rect 47 51 52 53
rect 16 39 21 41
rect 20 35 21 39
rect 16 33 21 35
rect 23 39 29 41
rect 23 35 24 39
rect 28 35 29 39
rect 23 33 29 35
rect 31 39 36 41
rect 31 35 32 39
rect 31 33 36 35
rect 40 39 45 41
rect 44 35 45 39
rect 40 33 45 35
rect 47 39 52 41
rect 47 35 48 39
rect 47 33 52 35
<< ndcontact >>
rect 16 173 20 177
rect 24 173 28 177
rect 32 173 36 177
rect 40 175 44 179
rect 48 175 52 179
rect 16 99 20 103
rect 24 99 28 103
rect 32 99 36 103
rect 40 97 44 101
rect 48 97 52 101
rect 7 83 11 87
rect 16 79 20 87
rect 24 81 28 85
rect 32 81 36 85
rect 40 83 44 87
rect 48 83 52 87
rect 16 7 20 11
rect 24 7 28 11
rect 32 7 36 11
rect 40 5 44 9
rect 48 5 52 9
<< pdcontact >>
rect 16 145 20 149
rect 24 145 28 149
rect 32 145 36 149
rect 40 145 44 149
rect 48 145 52 149
rect 16 127 20 131
rect 24 127 28 131
rect 32 127 36 131
rect 40 127 44 131
rect 48 127 52 131
rect 7 51 11 55
rect 16 51 20 55
rect 24 53 28 57
rect 32 53 36 57
rect 40 53 44 57
rect 48 53 52 57
rect 16 35 20 39
rect 24 35 28 39
rect 32 35 36 39
rect 40 35 44 39
rect 48 35 52 39
<< psubstratepcontact >>
rect 40 167 44 171
rect 40 105 44 109
rect 40 75 44 79
rect 40 13 44 17
<< nsubstratencontact >>
rect 56 145 60 149
rect 56 127 60 131
rect 56 53 60 57
rect 56 35 60 39
<< polysilicon >>
rect 21 179 23 181
rect 29 179 31 181
rect 45 179 47 181
rect 21 151 23 171
rect 29 166 31 171
rect 30 162 31 166
rect 29 151 31 162
rect 45 151 47 175
rect 21 141 23 143
rect 29 141 31 143
rect 45 141 47 143
rect 21 133 23 135
rect 29 133 31 135
rect 45 133 47 135
rect 21 105 23 125
rect 29 114 31 125
rect 30 110 31 114
rect 29 105 31 110
rect 45 101 47 125
rect 21 95 23 97
rect 29 95 31 97
rect 45 95 47 97
rect 12 87 14 89
rect 21 87 23 89
rect 29 87 31 89
rect 45 87 47 89
rect 12 59 14 83
rect 21 59 23 79
rect 29 76 31 79
rect 30 72 31 76
rect 29 59 31 72
rect 45 59 47 83
rect 12 49 14 51
rect 21 49 23 51
rect 29 49 31 51
rect 45 49 47 51
rect 21 41 23 43
rect 29 41 31 43
rect 45 41 47 43
rect 21 13 23 33
rect 29 22 31 33
rect 30 18 31 22
rect 29 13 31 18
rect 45 9 47 33
rect 21 3 23 5
rect 29 3 31 5
rect 45 3 47 5
<< polycontact >>
rect 17 154 21 158
rect 26 162 30 166
rect 41 159 45 163
rect 17 118 21 122
rect 26 110 30 114
rect 41 113 45 117
rect 8 66 12 70
rect 17 62 21 66
rect 26 72 30 76
rect 41 67 45 71
rect 17 26 21 30
rect 26 18 30 22
rect 41 21 45 25
<< metal1 >>
rect 0 182 64 186
rect 16 177 20 182
rect 40 179 44 182
rect 0 162 26 165
rect 33 162 36 173
rect 40 171 44 175
rect 52 175 55 179
rect 59 175 64 179
rect 33 159 41 162
rect 33 157 36 159
rect 24 154 36 157
rect 24 149 28 154
rect 40 149 44 151
rect 16 140 20 145
rect 32 140 36 145
rect 40 140 44 145
rect 48 149 52 175
rect 48 143 52 145
rect 56 140 60 145
rect 0 136 64 140
rect 16 131 20 136
rect 32 131 36 136
rect 40 131 44 136
rect 24 122 28 127
rect 40 125 44 127
rect 48 131 52 133
rect 56 131 60 136
rect 24 119 36 122
rect 33 117 36 119
rect 33 114 41 117
rect 0 110 26 113
rect 33 103 36 114
rect 40 101 44 105
rect 16 94 20 99
rect 48 101 52 127
rect 52 97 55 101
rect 59 97 64 101
rect 40 94 44 97
rect 0 90 64 94
rect 16 87 20 90
rect 40 87 44 90
rect 0 73 26 76
rect 33 70 36 81
rect 40 79 44 83
rect 52 83 55 87
rect 59 83 64 87
rect 0 66 8 68
rect 0 65 12 66
rect 33 67 41 70
rect 33 65 36 67
rect 24 62 36 65
rect 24 57 28 62
rect 40 57 44 59
rect 16 48 20 51
rect 32 48 36 53
rect 40 48 44 53
rect 48 57 52 83
rect 48 51 52 53
rect 56 48 60 53
rect 0 44 64 48
rect 16 39 20 44
rect 32 39 36 44
rect 40 39 44 44
rect 24 30 28 35
rect 40 33 44 35
rect 48 39 52 41
rect 56 39 60 44
rect 24 27 36 30
rect 33 25 36 27
rect 33 22 41 25
rect 0 19 26 22
rect 33 11 36 22
rect 40 9 44 13
rect 16 2 20 7
rect 48 9 52 35
rect 52 5 55 9
rect 59 5 64 9
rect 40 2 44 5
rect 0 -2 64 2
<< m2contact >>
rect 55 175 59 179
rect 13 154 17 158
rect 13 118 17 122
rect 55 97 59 101
rect 7 79 11 83
rect 55 83 59 87
rect 17 66 21 70
rect 7 55 11 59
rect 13 26 17 30
rect 55 5 59 9
<< metal2 >>
rect 13 122 17 154
rect 13 83 17 118
rect 11 79 17 83
rect 13 59 17 79
rect 11 55 17 59
rect 13 30 17 55
<< m3contact >>
rect 59 175 63 179
rect 59 97 63 101
rect 59 83 63 87
rect 59 5 63 9
<< metal3 >>
rect 58 179 64 180
rect 58 175 59 179
rect 63 175 64 179
rect 58 174 64 175
rect 58 101 64 102
rect 58 97 59 101
rect 63 97 64 101
rect 58 96 64 97
rect 58 87 64 88
rect 58 83 59 87
rect 63 83 64 87
rect 58 82 64 83
rect 58 9 64 10
rect 58 5 59 9
rect 63 5 64 9
rect 58 4 64 5
<< m3p >>
rect 0 0 64 184
<< labels >>
rlabel metal1 64 5 64 5 7 out0
rlabel metal1 64 84 64 84 1 out1
rlabel metal1 64 97 64 97 7 out2
rlabel metal1 64 175 64 175 7 out3
rlabel metal1 0 162 0 162 3 in3
rlabel metal1 0 184 0 184 2 gnd
rlabel metal1 0 138 0 138 2 vdd
rlabel metal1 0 110 0 110 3 in2
rlabel metal1 0 46 0 46 2 vdd
rlabel metal1 0 19 0 19 3 in0
rlabel metal1 0 0 0 0 6 gnd
rlabel metal1 0 92 0 92 4 gnd
rlabel metal1 0 73 0 73 3 in1
rlabel metal1 0 65 0 65 3 en
<< end >>
