magic
tech scmos
timestamp 1565708499
<< nwell >>
rect 0 -2 25 40
<< pwell >>
rect 25 -2 44 40
<< ntransistor >>
rect 31 18 35 20
rect 31 10 35 12
<< ptransistor >>
rect 11 18 19 20
rect 11 10 19 12
<< ndiffusion >>
rect 31 20 35 21
rect 31 17 35 18
rect 31 12 35 13
rect 31 9 35 10
<< pdiffusion >>
rect 11 21 13 25
rect 17 21 19 25
rect 11 20 19 21
rect 11 12 19 18
rect 11 9 19 10
rect 11 5 13 9
rect 17 5 19 9
<< ndcontact >>
rect 31 21 35 25
rect 31 13 35 17
rect 31 5 35 9
<< pdcontact >>
rect 13 21 17 25
rect 13 5 17 9
<< psubstratepcontact >>
rect 31 29 35 33
<< nsubstratencontact >>
rect 13 29 17 33
<< polysilicon >>
rect 10 18 11 20
rect 19 18 31 20
rect 35 18 39 20
rect 10 10 11 12
rect 19 10 31 12
rect 35 10 39 12
<< polycontact >>
rect 6 16 10 20
rect 6 8 10 12
<< metal1 >>
rect 0 36 44 40
rect 13 33 17 36
rect 13 25 17 29
rect 0 21 10 24
rect 27 25 31 33
rect 6 20 10 21
rect 38 17 44 20
rect 21 13 31 17
rect 35 14 41 17
rect 0 9 6 12
rect 21 9 24 13
rect 17 5 24 9
rect 27 2 31 5
rect 0 -2 44 2
<< m2contact >>
rect 27 21 31 25
rect 27 5 31 9
<< metal2 >>
rect 27 9 31 21
<< m3p >>
rect 0 0 44 38
<< labels >>
rlabel metal1 44 17 44 17 7 Z
rlabel metal1 0 9 0 9 3 B
rlabel metal1 0 21 0 21 1 A
rlabel metal1 0 38 0 38 1 vdd
rlabel metal1 0 0 0 0 1 gnd
<< end >>
