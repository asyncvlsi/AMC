magic
tech scmos
timestamp 1553263517
<< nwell >>
rect 0 -2 23 40
<< pwell >>
rect 23 -2 43 40
<< ntransistor >>
rect 29 26 37 28
rect 29 18 37 20
<< ptransistor >>
rect 9 26 17 28
rect 9 18 17 20
<< ndiffusion >>
rect 29 29 31 33
rect 35 29 37 33
rect 29 28 37 29
rect 29 20 37 26
rect 29 14 37 18
rect 29 10 31 14
rect 35 10 37 14
<< pdiffusion >>
rect 9 29 11 33
rect 15 29 17 33
rect 9 28 17 29
rect 9 25 17 26
rect 9 21 11 25
rect 15 21 17 25
rect 9 20 17 21
rect 9 17 17 18
rect 9 13 11 17
rect 15 13 17 17
<< ndcontact >>
rect 31 29 35 33
rect 31 10 35 14
<< pdcontact >>
rect 11 29 15 33
rect 11 21 15 25
rect 11 13 15 17
<< psubstratepcontact >>
rect 31 2 35 6
<< nsubstratencontact >>
rect 15 5 19 9
<< polysilicon >>
rect 8 26 9 28
rect 17 26 29 28
rect 37 26 39 28
rect 8 18 9 20
rect 17 18 29 20
rect 37 18 39 20
<< polycontact >>
rect 4 24 8 28
rect 4 16 8 20
<< metal1 >>
rect 0 36 15 40
rect 19 36 43 40
rect 0 24 4 27
rect 31 25 35 29
rect 15 21 35 25
rect 30 20 35 21
rect 0 16 4 17
rect 30 17 43 20
rect 0 14 8 16
rect 15 9 19 13
rect 31 6 35 10
rect 0 -2 43 2
<< m2contact >>
rect 15 36 19 40
rect 15 29 19 33
rect 15 13 19 17
<< metal2 >>
rect 15 33 19 36
rect 15 17 19 29
<< m3p >>
rect 0 0 43 38
<< labels >>
rlabel metal1 0 38 0 38 4 vdd
rlabel metal1 0 0 0 0 2 gnd
rlabel metal1 0 24 0 24 1 B
rlabel metal1 43 17 43 17 7 Z
rlabel metal1 0 14 0 14 1 A
<< end >>
