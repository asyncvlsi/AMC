magic
tech scmos
timestamp 1553355638
<< nwell >>
rect -1 -2 24 40
<< pwell >>
rect 24 -2 49 40
<< ntransistor >>
rect 35 26 43 28
rect 35 18 43 20
rect 35 10 43 12
<< ptransistor >>
rect 10 26 18 28
rect 10 18 18 20
rect 10 10 18 12
<< ndiffusion >>
rect 35 29 37 33
rect 41 29 43 33
rect 35 28 43 29
rect 35 20 43 26
rect 35 12 43 18
rect 35 9 43 10
rect 35 5 37 9
rect 41 5 43 9
<< pdiffusion >>
rect 10 29 12 33
rect 16 29 18 33
rect 10 28 18 29
rect 10 25 18 26
rect 10 21 12 25
rect 16 21 18 25
rect 10 20 18 21
rect 10 17 18 18
rect 10 13 12 17
rect 16 13 18 17
rect 10 12 18 13
rect 10 9 18 10
rect 10 5 12 9
rect 16 5 18 9
<< ndcontact >>
rect 37 29 41 33
rect 37 5 41 9
<< pdcontact >>
rect 12 29 16 33
rect 12 21 16 25
rect 12 13 16 17
rect 12 5 16 9
<< psubstratepcontact >>
rect 27 5 31 9
<< nsubstratencontact >>
rect 2 31 6 35
<< polysilicon >>
rect 8 26 10 28
rect 18 26 35 28
rect 43 26 45 28
rect 8 18 10 20
rect 18 18 35 20
rect 43 18 45 20
rect 8 10 10 12
rect 18 10 35 12
rect 43 10 45 12
<< polycontact >>
rect 4 24 8 28
rect 4 16 8 20
rect 4 8 8 12
<< metal1 >>
rect 0 36 16 40
rect 20 36 49 40
rect 2 35 6 36
rect 16 29 26 33
rect 0 24 4 27
rect 23 21 26 29
rect 37 21 41 29
rect 23 20 41 21
rect 0 16 4 19
rect 23 17 49 20
rect 16 13 26 17
rect 0 8 4 11
rect 27 2 31 5
rect 37 2 41 5
rect 0 -2 49 2
<< m2contact >>
rect 16 36 20 40
rect 16 21 20 25
rect 16 5 20 9
<< metal2 >>
rect 16 25 20 36
rect 16 9 20 21
<< m3p >>
rect 0 0 49 38
<< labels >>
rlabel metal1 0 0 0 0 1 gnd
rlabel metal1 0 38 0 38 1 vdd
rlabel metal1 0 8 0 8 1 A
rlabel metal1 0 16 0 16 1 B
rlabel metal1 0 24 0 24 1 C
rlabel metal1 49 17 49 17 7 Z
<< end >>
